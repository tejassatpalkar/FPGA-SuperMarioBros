/*

struct {
	logic [9:0]  x, y,
	enum logic [2:0] {BLOCK, MARIO, GROUND, MUSHROOM} sprite_type,
	int width, height,
} sprite_position
*/